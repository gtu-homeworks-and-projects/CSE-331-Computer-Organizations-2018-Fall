module shifter_32 (out, in1, in2, shiftMode, logical);
input [31:0] in1;
input [4:0] in2;
input shiftMode, logical;
output [31:0] out;

wire [31:0] out1, out2, out3, out4;
wire [1:0] mode1, mode2, mode3, mode4, mode5;
wire leftMostBit, notShiftMode, arithmeticLeftMost;

not (notShiftMode, shiftMode);
and determine_left_most(arithmeticLeftMost, in1[31], notShiftMode);
mux_2x1 aOrL(leftMostBit, arithmeticLeftMost, 1'b0, logical);
buf (mode1[0], shiftMode);
buf (mode2[0], shiftMode);
buf (mode3[0], shiftMode);
buf (mode4[0], shiftMode);
buf (mode5[0], shiftMode);

buf (mode1[1], in2[0]);
mux_4x1 firstMux1(out1[0], in1[0], in1[0], in1[1], 1'b0, mode1),
	firstMux2(out1[1], in1[1], in1[1], in1[2], in1[0], mode1),
	firstMux3(out1[2], in1[2], in1[2], in1[3], in1[1], mode1),
	firstMux4(out1[3], in1[3], in1[3], in1[4], in1[2], mode1),
	firstMux5(out1[4], in1[4], in1[4], in1[5], in1[3], mode1),
	firstMux6(out1[5], in1[5], in1[5], in1[6], in1[4], mode1),
	firstMux7(out1[6], in1[6], in1[6], in1[7], in1[5], mode1),
	firstMux8(out1[7], in1[7], in1[7], in1[8], in1[6], mode1),
	firstMux9(out1[8], in1[8], in1[8], in1[9], in1[7], mode1),
	firstMux10(out1[9], in1[9], in1[9], in1[10], in1[8], mode1),
	firstMux11(out1[10], in1[10], in1[10], in1[11], in1[9], mode1),
	firstMux12(out1[11], in1[11], in1[11], in1[12], in1[10], mode1),
	firstMux13(out1[12], in1[12], in1[12], in1[13], in1[11], mode1),
	firstMux14(out1[13], in1[13], in1[13], in1[14], in1[12], mode1),
	firstMux15(out1[14], in1[14], in1[14], in1[15], in1[13], mode1),
	firstMux16(out1[15], in1[15], in1[15], in1[16], in1[14], mode1),
	firstMux17(out1[16], in1[16], in1[16], in1[17], in1[15], mode1),
	firstMux18(out1[17], in1[17], in1[17], in1[18], in1[16], mode1),
	firstMux19(out1[18], in1[18], in1[18], in1[19], in1[17], mode1),
	firstMux20(out1[19], in1[19], in1[19], in1[20], in1[18], mode1),
	firstMux21(out1[20], in1[20], in1[20], in1[21], in1[19], mode1),
	firstMux22(out1[21], in1[21], in1[21], in1[22], in1[20], mode1),
	firstMux23(out1[22], in1[22], in1[22], in1[23], in1[21], mode1),
	firstMux24(out1[23], in1[23], in1[23], in1[24], in1[22], mode1),
	firstMux25(out1[24], in1[24], in1[24], in1[25], in1[23], mode1),
	firstMux26(out1[25], in1[25], in1[25], in1[26], in1[24], mode1),
	firstMux27(out1[26], in1[26], in1[26], in1[27], in1[25], mode1),
	firstMux28(out1[27], in1[27], in1[27], in1[28], in1[26], mode1),
	firstMux29(out1[28], in1[28], in1[28], in1[29], in1[27], mode1),
	firstMux30(out1[29], in1[29], in1[29], in1[30], in1[28], mode1),
	firstMux31(out1[30], in1[30], in1[30], in1[31], in1[29], mode1),
	firstMux32(out1[31], in1[31], in1[31], leftMostBit, in1[30], mode1);

buf (mode2[1], in2[1]);
mux_4x1 secondMux1(out2[0], out1[0], out1[0], out1[2], 1'b0, mode2),
	secondMux2(out2[1], out1[1], out1[1], out1[3], 1'b0, mode2),
	secondMux3(out2[2], out1[2], out1[2], out1[4], out1[0], mode2),
	secondMux4(out2[3], out1[3], out1[3], out1[5], out1[1], mode2),
	secondMux5(out2[4], out1[4], out1[4], out1[6], out1[2], mode2),
	secondMux6(out2[5], out1[5], out1[5], out1[7], out1[3], mode2),
	secondMux7(out2[6], out1[6], out1[6], out1[8], out1[4], mode2),
	secondMux8(out2[7], out1[7], out1[7], out1[9], out1[5], mode2),
	secondMux9(out2[8], out1[8], out1[8], out1[10], out1[6], mode2),
	secondMux10(out2[9], out1[9], out1[9], out1[11], out1[7], mode2),
	secondMux11(out2[10], out1[10], out1[10], out1[12], out1[8], mode2),
	secondMux12(out2[11], out1[11], out1[11], out1[13], out1[9], mode2),
	secondMux13(out2[12], out1[12], out1[12], out1[14], out1[10], mode2),
	secondMux14(out2[13], out1[13], out1[13], out1[15], out1[11], mode2),
	secondMux15(out2[14], out1[14], out1[14], out1[16], out1[12], mode2),
	secondMux16(out2[15], out1[15], out1[15], out1[17], out1[13], mode2),
	secondMux17(out2[16], out1[16], out1[16], out1[18], out1[14], mode2),
	secondMux18(out2[17], out1[17], out1[17], out1[19], out1[15], mode2),
	secondMux19(out2[18], out1[18], out1[18], out1[20], out1[16], mode2),
	secondMux20(out2[19], out1[19], out1[19], out1[21], out1[17], mode2),
	secondMux21(out2[20], out1[20], out1[20], out1[22], out1[18], mode2),
	secondMux22(out2[21], out1[21], out1[21], out1[23], out1[19], mode2),
	secondMux23(out2[22], out1[22], out1[22], out1[24], out1[20], mode2),
	secondMux24(out2[23], out1[23], out1[23], out1[25], out1[21], mode2),
	secondMux25(out2[24], out1[24], out1[24], out1[26], out1[22], mode2),
	secondMux26(out2[25], out1[25], out1[25], out1[27], out1[23], mode2),
	secondMux27(out2[26], out1[26], out1[26], out1[28], out1[24], mode2),
	secondMux28(out2[27], out1[27], out1[27], out1[29], out1[25], mode2),
	secondMux29(out2[28], out1[28], out1[28], out1[30], out1[26], mode2),
	secondMux30(out2[29], out1[29], out1[29], out1[31], out1[27], mode2),
	secondMux31(out2[30], out1[30], out1[30], leftMostBit, out1[28], mode2),
	secondMux32(out2[31], out1[31], out1[31], leftMostBit, out1[29], mode2);

buf (mode3[1], in2[2]);
mux_4x1 thirdMux1(out3[0], out2[0], out2[0], out2[4], 1'b0, mode3),
	thirdMux2(out3[1], out2[1], out2[1], out2[5], 1'b0, mode3),
	thirdMux3(out3[2], out2[2], out2[2], out2[6], 1'b0, mode3),
	thirdMux4(out3[3], out2[3], out2[3], out2[7], 1'b0, mode3),
	thirdMux5(out3[4], out2[4], out2[4], out2[8], out2[0], mode3),
	thirdMux6(out3[5], out2[5], out2[5], out2[9], out2[1], mode3),
	thirdMux7(out3[6], out2[6], out2[6], out2[10], out2[2], mode3),
	thirdMux8(out3[7], out2[7], out2[7], out2[11], out2[3], mode3),
	thirdMux9(out3[8], out2[8], out2[8], out2[12], out2[4], mode3),
	thirdMux10(out3[9], out2[9], out2[9], out2[13], out2[5], mode3),
	thirdMux11(out3[10], out2[10], out2[10], out2[14], out2[6], mode3),
	thirdMux12(out3[11], out2[11], out2[11], out2[15], out2[7], mode3),
	thirdMux13(out3[12], out2[12], out2[12], out2[16], out2[8], mode3),
	thirdMux14(out3[13], out2[13], out2[13], out2[17], out2[9], mode3),
	thirdMux15(out3[14], out2[14], out2[14], out2[18], out2[10], mode3),
	thirdMux16(out3[15], out2[15], out2[15], out2[19], out2[11], mode3),
	thirdMux17(out3[16], out2[16], out2[16], out2[20], out2[12], mode3),
	thirdMux18(out3[17], out2[17], out2[17], out2[21], out2[13], mode3),
	thirdMux19(out3[18], out2[18], out2[18], out2[22], out2[14], mode3),
	thirdMux20(out3[19], out2[19], out2[19], out2[23], out2[15], mode3),
	thirdMux21(out3[20], out2[20], out2[20], out2[24], out2[16], mode3),
	thirdMux22(out3[21], out2[21], out2[21], out2[25], out2[17], mode3),
	thirdMux23(out3[22], out2[22], out2[22], out2[26], out2[18], mode3),
	thirdMux24(out3[23], out2[23], out2[23], out2[27], out2[19], mode3),
	thirdMux25(out3[24], out2[24], out2[24], out2[28], out2[20], mode3),
	thirdMux26(out3[25], out2[25], out2[25], out2[29], out2[21], mode3),
	thirdMux27(out3[26], out2[26], out2[26], out2[30], out2[22], mode3),
	thirdMux28(out3[27], out2[27], out2[27], out2[31], out2[23], mode3),
	thirdMux29(out3[28], out2[28], out2[28], leftMostBit, out2[24], mode3),
	thirdMux30(out3[29], out2[29], out2[29], leftMostBit, out2[25], mode3),
	thirdMux31(out3[30], out2[30], out2[30], leftMostBit, out2[26], mode3),
	thirdMux32(out3[31], out2[31], out2[31], leftMostBit, out2[27], mode3);
	
buf (mode4[1], in2[3]);
mux_4x1 fourthMux1(out4[0], out3[0], out3[0], out3[8], 1'b0, mode4),
	fourthMux2(out4[1], out3[1], out3[1], out3[9], 1'b0, mode4),
	fourthMux3(out4[2], out3[2], out3[2], out3[10], 1'b0, mode4),
	fourthMux4(out4[3], out3[3], out3[3], out3[11], 1'b0, mode4),
	fourthMux5(out4[4], out3[4], out3[4], out3[12], 1'b0, mode4),
	fourthMux6(out4[5], out3[5], out3[5], out3[13], 1'b0, mode4),
	fourthMux7(out4[6], out3[6], out3[6], out3[14], 1'b0, mode4),
	fourthMux8(out4[7], out3[7], out3[7], out3[15], 1'b0, mode4),
	fourthMux9(out4[8], out3[8], out3[8], out3[16], out3[0], mode4),
	fourthMux10(out4[9], out3[9], out3[9], out3[17], out3[1], mode4),
	fourthMux11(out4[10], out3[10], out3[10], out3[18], out3[2], mode4),
	fourthMux12(out4[11], out3[11], out3[11], out3[19], out3[3], mode4),
	fourthMux13(out4[12], out3[12], out3[12], out3[20], out3[4], mode4),
	fourthMux14(out4[13], out3[13], out3[13], out3[21], out3[5], mode4),
	fourthMux15(out4[14], out3[14], out3[14], out3[22], out3[6], mode4),
	fourthMux16(out4[15], out3[15], out3[15], out3[23], out3[7], mode4),
	fourthMux17(out4[16], out3[16], out3[16], out3[24], out3[8], mode4),
	fourthMux18(out4[17], out3[17], out3[17], out3[25], out3[9], mode4),
	fourthMux19(out4[18], out3[18], out3[18], out3[26], out3[10], mode4),
	fourthMux20(out4[19], out3[19], out3[19], out3[27], out3[11], mode4),
	fourthMux21(out4[20], out3[20], out3[20], out3[28], out3[12], mode4),
	fourthMux22(out4[21], out3[21], out3[21], out3[29], out3[13], mode4),
	fourthMux23(out4[22], out3[22], out3[22], out3[30], out3[14], mode4),
	fourthMux24(out4[23], out3[23], out3[23], out3[31], out3[15], mode4),
	fourthMux25(out4[24], out3[24], out3[24], leftMostBit, out3[16], mode4),
	fourthMux26(out4[25], out3[25], out3[25], leftMostBit, out3[17], mode4),
	fourthMux27(out4[26], out3[26], out3[26], leftMostBit, out3[18], mode4),
	fourthMux28(out4[27], out3[27], out3[27], leftMostBit, out3[19], mode4),
	fourthMux29(out4[28], out3[28], out3[28], leftMostBit, out3[20], mode4),
	fourthMux30(out4[29], out3[29], out3[29], leftMostBit, out3[21], mode4),
	fourthMux31(out4[30], out3[30], out3[30], leftMostBit, out3[22], mode4),
	fourthMux32(out4[31], out3[31], out3[31], leftMostBit, out3[23], mode4);
		
buf (mode5[1], in2[4]);
mux_4x1 fifthMux1(out[0], out4[0], out4[0], out4[16], 1'b0, mode5),
	fifthMux2(out[1], out4[1], out4[1], out4[17], 1'b0, mode5),
	fifthMux3(out[2], out4[2], out4[2], out4[18], 1'b0, mode5),
	fifthMux4(out[3], out4[3], out4[3], out4[19], 1'b0, mode5),
	fifthMux5(out[4], out4[4], out4[4], out4[20], 1'b0, mode5),
	fifthMux6(out[5], out4[5], out4[5], out4[21], 1'b0, mode5),
	fifthMux7(out[6], out4[6], out4[6], out4[22], 1'b0, mode5),
	fifthMux8(out[7], out4[7], out4[7], out4[23], 1'b0, mode5),
	fifthMux9(out[8], out4[8], out4[8], out4[24], 1'b0, mode5),
	fifthMux10(out[9], out4[9], out4[9], out4[25], 1'b0, mode5),
	fifthMux11(out[10], out4[10], out4[10], out4[26], 1'b0, mode5),
	fifthMux12(out[11], out4[11], out4[11], out4[27], 1'b0, mode5),
	fifthMux13(out[12], out4[12], out4[12], out4[28], 1'b0, mode5),
	fifthMux14(out[13], out4[13], out4[13], out4[29], 1'b0, mode5),
	fifthMux15(out[14], out4[14], out4[14], out4[30], 1'b0, mode5),
	fifthMux16(out[15], out4[15], out4[15], out4[31], 1'b0, mode5),
	fifthMux17(out[16], out4[16], out4[16], leftMostBit, out4[0], mode5),
	fifthMux18(out[17], out4[17], out4[17], leftMostBit, out4[1], mode5),
	fifthMux19(out[18], out4[18], out4[18], leftMostBit, out4[2], mode5),
	fifthMux20(out[19], out4[19], out4[19], leftMostBit, out4[3], mode5),
	fifthMux21(out[20], out4[20], out4[20], leftMostBit, out4[4], mode5),
	fifthMux22(out[21], out4[21], out4[21], leftMostBit, out4[5], mode5),
	fifthMux23(out[22], out4[22], out4[22], leftMostBit, out4[6], mode5),
	fifthMux24(out[23], out4[23], out4[23], leftMostBit, out4[7], mode5),
	fifthMux25(out[24], out4[24], out4[24], leftMostBit, out4[8], mode5),
	fifthMux26(out[25], out4[25], out4[25], leftMostBit, out4[9], mode5),
	fifthMux27(out[26], out4[26], out4[26], leftMostBit, out4[10], mode5),
	fifthMux28(out[27], out4[27], out4[27], leftMostBit, out4[11], mode5),
	fifthMux29(out[28], out4[28], out4[28], leftMostBit, out4[12], mode5),
	fifthMux30(out[29], out4[29], out4[29], leftMostBit, out4[13], mode5),
	fifthMux31(out[30], out4[30], out4[30], leftMostBit, out4[14], mode5),
	fifthMux32(out[31], out4[31], out4[31], leftMostBit, out4[15], mode5);

endmodule