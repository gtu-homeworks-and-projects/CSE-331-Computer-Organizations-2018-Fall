`define DELAY 10

module alu32_testbench();
reg [31:0] A,B;
reg [2:0] S;
wire [31:0] R;
alu32 alu(R, A, B, S);

initial begin
// AND
S = 3'b000; 
A = 32'b01111011111111111111111111111110;
B = 32'b11111111111111111100001111111111;
#`DELAY;
A = 32'b01111011111111111111100011111110;
B = 32'b11111111100011111100001111111111;
#`DELAY;
A = 32'b01111011111110000011111111111110;
B = 32'b00100011100011111100001111111111;
#`DELAY;

// OR
S = 3'b001;
A = 32'b01111011111110000011111111111110;
B = 32'b11111111100011111100001111100011;
#`DELAY;
A = 32'b01111011111111000000000000000110;
B = 32'b11111111100011111100001111111111;
#`DELAY;
A = 32'b01111011111110000011111111111110;
B = 32'b11111111100011111100001111111111;
#`DELAY;

// Addition
S = 3'b010;
A = 32'b00000000000000000000000000000010;
B = 4;
#`DELAY;
A = 12;
B = 25;
#`DELAY;
A = 8692468;
B = 307532;
#`DELAY;

// XOR
S = 3'b011;
A = 32'b01010101010101010101010101010101;
B = 32'b10101010101010101010101010101010;
#`DELAY;
A = 32'b00011011100111111110000111001010;
B = 32'b11001101100000001111110000000111;
#`DELAY;
A = 32'b01101110111111111110000111111111;
B = 32'b01111111111111111111111111111111;
#`DELAY;

// Subtraction
S = 3'b100;
A = 32'b00000000000000000000000000000110;
B = 4;
#`DELAY;
A = 25;
B = 12;
#`DELAY;
A = 8692468;
B = 692468;
#`DELAY;

// Arithmetic Right Shift
S = 3'b101;
A = 32'b00000000000000000000000000001000;
B = 32'b00000000000000000000000000000001;
#`DELAY;
A = 32'b11111111111111111110000011111100;
B = 32'b00000000000000000000000000011111;
#`DELAY;
A = 32'b11111111100000000011110000000000;
B = 32'b00000000000000000000000000000011;
#`DELAY;

// Left Shift
S = 3'b110;
A = 32'b00000000000000000000000000001000;
B = 32'b00000000000000000000000000000001;
#`DELAY;
A = 32'b11111111111111111110000011111101;
B = 32'b00000000000000000000000000011110;
#`DELAY;
A = 32'b10000000000000000000000000000000;
B = 32'b00000000000000000000000000000011;
#`DELAY;

// NOR
S = 3'b111;
A = 32'b11111100000000000000000000001000;
B = 32'b00000000111111111100000000000001;
#`DELAY;
A = 32'b11111111111111111110010011111101;
B = 32'b00000000000000011111100000011110;
#`DELAY;
A = 32'b10000000000000000000000001000000;
B = 32'b00000000010000000000000000000011;
#`DELAY;
end

initial begin
$monitor("time = %2d, A = %32b, B=%32b, R=%32b, S=%3b", $time, A, B, R, S);
end

endmodule