module not_32 (out, in);
input [31:0] in;
output [31:0] out;

not not1(out[0], in[0]),
	not2(out[1], in[1]),
	not3(out[2], in[2]),
	not4(out[3], in[3]),
	not5(out[4], in[4]),
	not6(out[5], in[5]),
	not7(out[6], in[6]),
	not8(out[7], in[7]),
	not9(out[8], in[8]),
	not10(out[9], in[9]),
	not11(out[10], in[10]),
	not12(out[11], in[11]),
	not13(out[12], in[12]),
	not14(out[13], in[13]),
	not15(out[14], in[14]),
	not16(out[15], in[15]),
	not17(out[16], in[16]),
	not18(out[17], in[17]),
	not19(out[18], in[18]),
	not20(out[19], in[19]),
	not21(out[20], in[20]),
	not22(out[21], in[21]),
	not23(out[22], in[22]),
	not24(out[23], in[23]),
	not25(out[24], in[24]),
	not26(out[25], in[25]),
	not27(out[26], in[26]),
	not28(out[27], in[27]),
	not29(out[28], in[28]),
	not30(out[29], in[29]),
	not31(out[30], in[30]),
	not32(out[31], in[31]);
	
endmodule